package fifo_env_pkg;

import uvm_pkg::*;
import fifo_agent_pkg::*;

`include "uvm_macros.svh"
`include "fifo_env.sv"

endpackage: fifo_env_pkg