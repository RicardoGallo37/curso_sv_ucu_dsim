// Interface definitions for counter  
interface cnt_if #(parameter WIDTH = 4) (input bit clk);
  logic             rstn;
  logic             load_en;
  logic [WIDTH-1:0] load;
  logic [WIDTH-1:0] count;
  logic             down;
  logic             rollover;
endinterface
