package tests_pkg;

import uvm_pkg::*;
import fifo_env_pkg::*;
import fifo_agent_pkg::*;

`include "uvm_macros.svh"
`include "fifo_test.sv"

endpackage: tests_pkg