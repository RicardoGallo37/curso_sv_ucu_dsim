package fifo_agent_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

`include "fifo_agent_config.sv"
`include "fifo_transaction.sv"
`include "fifo_sequence.sv"
`include "fifo_driver.sv"
`include "fifo_monitor.sv"
`include "fifo_sequencer.sv"
`include "fifo_agent.sv"

endpackage