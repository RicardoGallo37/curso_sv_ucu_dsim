package tests_pkg;

import uvm_pkg::*;
import fifo_env_pkg::*;
import fifo_agent_pkg::*;

`include "uvm_macros.svh"
`include "fifo_test.sv"

//LAB: include another test that is a child of the fifo_test to change the config. Add the command to the makefile

endpackage: tests_pkg