
module fifo_top (fifo_ports ports, fifo_monitor_ports mports);

  import fifo_driver_pkg::*;

   //generate the driver component here
  ???

  initial begin
    //start the driver (use the function go)
    ???;
  end

//endprogram
endmodule
