
package definitions_pkg;

  parameter VERSION = "Rydev DSim System Verilog Course";
endpackage
